/**
 * 1-bit register:
 * If load[t] == 1 then out[t+1] = in[t]
 *    else out does not change (out[t+1] = out[t])
 */

`default_nettype none
module Bit(
	input wire clk,
	input wire in,
	input wire load,
	output wire out
);

// your implementation comes here:



endmodule
