/**
 * Adds two 16-bit values.
 * The most significant carry bit is ignored.
 * out = a + b (16 bit)
 */

`default_nettype none
module Add16(
	input wire [15:0] a,
	input wire [15:0] b,
	output wire [15:0] out
);
// your implementation comes here:


endmodule
